// TimerWithClock.v

// Generated using ACDS version 23.1 993

`timescale 1 ps / 1 ps
module TimerWithClock (
		input  wire [3:0] buttons_export,         //         buttons.export
		output wire       buzzer_export,          //          buzzer.export
		input  wire       clk_clk,                //             clk.clk
		output wire [9:0] leds_export,            //            leds.export
		output wire [6:0] sseg_hour_tens_export,  //  sseg_hour_tens.export
		output wire [6:0] sseg_hour_units_export, // sseg_hour_units.export
		output wire [6:0] sseg_min_units_export,  //  sseg_min_units.export
		output wire [6:0] sseg_mins_tens_export,  //  sseg_mins_tens.export
		output wire [6:0] sseg_sec_tens_export,   //   sseg_sec_tens.export
		output wire [6:0] sseg_sec_units_export,  //  sseg_sec_units.export
		input  wire       switch_export           //          switch.export
	);

	wire         timerwithclock_debug_reset_request_reset;                     // TimerWithClock:debug_reset_request -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire  [31:0] timerwithclock_data_master_readdata;                          // mm_interconnect_0:TimerWithClock_data_master_readdata -> TimerWithClock:d_readdata
	wire         timerwithclock_data_master_waitrequest;                       // mm_interconnect_0:TimerWithClock_data_master_waitrequest -> TimerWithClock:d_waitrequest
	wire         timerwithclock_data_master_debugaccess;                       // TimerWithClock:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:TimerWithClock_data_master_debugaccess
	wire  [13:0] timerwithclock_data_master_address;                           // TimerWithClock:d_address -> mm_interconnect_0:TimerWithClock_data_master_address
	wire   [3:0] timerwithclock_data_master_byteenable;                        // TimerWithClock:d_byteenable -> mm_interconnect_0:TimerWithClock_data_master_byteenable
	wire         timerwithclock_data_master_read;                              // TimerWithClock:d_read -> mm_interconnect_0:TimerWithClock_data_master_read
	wire         timerwithclock_data_master_write;                             // TimerWithClock:d_write -> mm_interconnect_0:TimerWithClock_data_master_write
	wire  [31:0] timerwithclock_data_master_writedata;                         // TimerWithClock:d_writedata -> mm_interconnect_0:TimerWithClock_data_master_writedata
	wire  [31:0] timerwithclock_instruction_master_readdata;                   // mm_interconnect_0:TimerWithClock_instruction_master_readdata -> TimerWithClock:i_readdata
	wire         timerwithclock_instruction_master_waitrequest;                // mm_interconnect_0:TimerWithClock_instruction_master_waitrequest -> TimerWithClock:i_waitrequest
	wire  [13:0] timerwithclock_instruction_master_address;                    // TimerWithClock:i_address -> mm_interconnect_0:TimerWithClock_instruction_master_address
	wire         timerwithclock_instruction_master_read;                       // TimerWithClock:i_read -> mm_interconnect_0:TimerWithClock_instruction_master_read
	wire         mm_interconnect_0_debug_avalon_jtag_slave_chipselect;         // mm_interconnect_0:DEBUG_avalon_jtag_slave_chipselect -> DEBUG:av_chipselect
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_readdata;           // DEBUG:av_readdata -> mm_interconnect_0:DEBUG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_debug_avalon_jtag_slave_waitrequest;        // DEBUG:av_waitrequest -> mm_interconnect_0:DEBUG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_debug_avalon_jtag_slave_address;            // mm_interconnect_0:DEBUG_avalon_jtag_slave_address -> DEBUG:av_address
	wire         mm_interconnect_0_debug_avalon_jtag_slave_read;               // mm_interconnect_0:DEBUG_avalon_jtag_slave_read -> DEBUG:av_read_n
	wire         mm_interconnect_0_debug_avalon_jtag_slave_write;              // mm_interconnect_0:DEBUG_avalon_jtag_slave_write -> DEBUG:av_write_n
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_writedata;          // mm_interconnect_0:DEBUG_avalon_jtag_slave_writedata -> DEBUG:av_writedata
	wire  [31:0] mm_interconnect_0_timerwithclock_debug_mem_slave_readdata;    // TimerWithClock:debug_mem_slave_readdata -> mm_interconnect_0:TimerWithClock_debug_mem_slave_readdata
	wire         mm_interconnect_0_timerwithclock_debug_mem_slave_waitrequest; // TimerWithClock:debug_mem_slave_waitrequest -> mm_interconnect_0:TimerWithClock_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_timerwithclock_debug_mem_slave_debugaccess; // mm_interconnect_0:TimerWithClock_debug_mem_slave_debugaccess -> TimerWithClock:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_timerwithclock_debug_mem_slave_address;     // mm_interconnect_0:TimerWithClock_debug_mem_slave_address -> TimerWithClock:debug_mem_slave_address
	wire         mm_interconnect_0_timerwithclock_debug_mem_slave_read;        // mm_interconnect_0:TimerWithClock_debug_mem_slave_read -> TimerWithClock:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_timerwithclock_debug_mem_slave_byteenable;  // mm_interconnect_0:TimerWithClock_debug_mem_slave_byteenable -> TimerWithClock:debug_mem_slave_byteenable
	wire         mm_interconnect_0_timerwithclock_debug_mem_slave_write;       // mm_interconnect_0:TimerWithClock_debug_mem_slave_write -> TimerWithClock:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_timerwithclock_debug_mem_slave_writedata;   // mm_interconnect_0:TimerWithClock_debug_mem_slave_writedata -> TimerWithClock:debug_mem_slave_writedata
	wire         mm_interconnect_0_sram_s1_chipselect;                         // mm_interconnect_0:SRAM_s1_chipselect -> SRAM:chipselect
	wire  [31:0] mm_interconnect_0_sram_s1_readdata;                           // SRAM:readdata -> mm_interconnect_0:SRAM_s1_readdata
	wire   [9:0] mm_interconnect_0_sram_s1_address;                            // mm_interconnect_0:SRAM_s1_address -> SRAM:address
	wire   [3:0] mm_interconnect_0_sram_s1_byteenable;                         // mm_interconnect_0:SRAM_s1_byteenable -> SRAM:byteenable
	wire         mm_interconnect_0_sram_s1_write;                              // mm_interconnect_0:SRAM_s1_write -> SRAM:write
	wire  [31:0] mm_interconnect_0_sram_s1_writedata;                          // mm_interconnect_0:SRAM_s1_writedata -> SRAM:writedata
	wire         mm_interconnect_0_sram_s1_clken;                              // mm_interconnect_0:SRAM_s1_clken -> SRAM:clken
	wire         mm_interconnect_0_leds_s1_chipselect;                         // mm_interconnect_0:LEDS_s1_chipselect -> LEDS:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                           // LEDS:readdata -> mm_interconnect_0:LEDS_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                            // mm_interconnect_0:LEDS_s1_address -> LEDS:address
	wire         mm_interconnect_0_leds_s1_write;                              // mm_interconnect_0:LEDS_s1_write -> LEDS:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                          // mm_interconnect_0:LEDS_s1_writedata -> LEDS:writedata
	wire         mm_interconnect_0_sseg_hour_units_s1_chipselect;              // mm_interconnect_0:SSEG_HOUR_UNITS_s1_chipselect -> SSEG_HOUR_UNITS:chipselect
	wire  [31:0] mm_interconnect_0_sseg_hour_units_s1_readdata;                // SSEG_HOUR_UNITS:readdata -> mm_interconnect_0:SSEG_HOUR_UNITS_s1_readdata
	wire   [1:0] mm_interconnect_0_sseg_hour_units_s1_address;                 // mm_interconnect_0:SSEG_HOUR_UNITS_s1_address -> SSEG_HOUR_UNITS:address
	wire         mm_interconnect_0_sseg_hour_units_s1_write;                   // mm_interconnect_0:SSEG_HOUR_UNITS_s1_write -> SSEG_HOUR_UNITS:write_n
	wire  [31:0] mm_interconnect_0_sseg_hour_units_s1_writedata;               // mm_interconnect_0:SSEG_HOUR_UNITS_s1_writedata -> SSEG_HOUR_UNITS:writedata
	wire         mm_interconnect_0_sseg_min_units_s1_chipselect;               // mm_interconnect_0:SSEG_MIN_UNITS_s1_chipselect -> SSEG_MIN_UNITS:chipselect
	wire  [31:0] mm_interconnect_0_sseg_min_units_s1_readdata;                 // SSEG_MIN_UNITS:readdata -> mm_interconnect_0:SSEG_MIN_UNITS_s1_readdata
	wire   [1:0] mm_interconnect_0_sseg_min_units_s1_address;                  // mm_interconnect_0:SSEG_MIN_UNITS_s1_address -> SSEG_MIN_UNITS:address
	wire         mm_interconnect_0_sseg_min_units_s1_write;                    // mm_interconnect_0:SSEG_MIN_UNITS_s1_write -> SSEG_MIN_UNITS:write_n
	wire  [31:0] mm_interconnect_0_sseg_min_units_s1_writedata;                // mm_interconnect_0:SSEG_MIN_UNITS_s1_writedata -> SSEG_MIN_UNITS:writedata
	wire         mm_interconnect_0_sseg_sec_units_s1_chipselect;               // mm_interconnect_0:SSEG_SEC_UNITS_s1_chipselect -> SSEG_SEC_UNITS:chipselect
	wire  [31:0] mm_interconnect_0_sseg_sec_units_s1_readdata;                 // SSEG_SEC_UNITS:readdata -> mm_interconnect_0:SSEG_SEC_UNITS_s1_readdata
	wire   [1:0] mm_interconnect_0_sseg_sec_units_s1_address;                  // mm_interconnect_0:SSEG_SEC_UNITS_s1_address -> SSEG_SEC_UNITS:address
	wire         mm_interconnect_0_sseg_sec_units_s1_write;                    // mm_interconnect_0:SSEG_SEC_UNITS_s1_write -> SSEG_SEC_UNITS:write_n
	wire  [31:0] mm_interconnect_0_sseg_sec_units_s1_writedata;                // mm_interconnect_0:SSEG_SEC_UNITS_s1_writedata -> SSEG_SEC_UNITS:writedata
	wire         mm_interconnect_0_sseg_mins_tens_s1_chipselect;               // mm_interconnect_0:SSEG_MINS_TENS_s1_chipselect -> SSEG_MINS_TENS:chipselect
	wire  [31:0] mm_interconnect_0_sseg_mins_tens_s1_readdata;                 // SSEG_MINS_TENS:readdata -> mm_interconnect_0:SSEG_MINS_TENS_s1_readdata
	wire   [1:0] mm_interconnect_0_sseg_mins_tens_s1_address;                  // mm_interconnect_0:SSEG_MINS_TENS_s1_address -> SSEG_MINS_TENS:address
	wire         mm_interconnect_0_sseg_mins_tens_s1_write;                    // mm_interconnect_0:SSEG_MINS_TENS_s1_write -> SSEG_MINS_TENS:write_n
	wire  [31:0] mm_interconnect_0_sseg_mins_tens_s1_writedata;                // mm_interconnect_0:SSEG_MINS_TENS_s1_writedata -> SSEG_MINS_TENS:writedata
	wire  [31:0] mm_interconnect_0_buttons_s1_readdata;                        // BUTTONS:readdata -> mm_interconnect_0:BUTTONS_s1_readdata
	wire   [1:0] mm_interconnect_0_buttons_s1_address;                         // mm_interconnect_0:BUTTONS_s1_address -> BUTTONS:address
	wire         mm_interconnect_0_timer_s1_chipselect;                        // mm_interconnect_0:TIMER_s1_chipselect -> TIMER:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                          // TIMER:readdata -> mm_interconnect_0:TIMER_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                           // mm_interconnect_0:TIMER_s1_address -> TIMER:address
	wire         mm_interconnect_0_timer_s1_write;                             // mm_interconnect_0:TIMER_s1_write -> TIMER:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                         // mm_interconnect_0:TIMER_s1_writedata -> TIMER:writedata
	wire         mm_interconnect_0_sseg_sec_tens_s1_chipselect;                // mm_interconnect_0:SSEG_SEC_TENS_s1_chipselect -> SSEG_SEC_TENS:chipselect
	wire  [31:0] mm_interconnect_0_sseg_sec_tens_s1_readdata;                  // SSEG_SEC_TENS:readdata -> mm_interconnect_0:SSEG_SEC_TENS_s1_readdata
	wire   [1:0] mm_interconnect_0_sseg_sec_tens_s1_address;                   // mm_interconnect_0:SSEG_SEC_TENS_s1_address -> SSEG_SEC_TENS:address
	wire         mm_interconnect_0_sseg_sec_tens_s1_write;                     // mm_interconnect_0:SSEG_SEC_TENS_s1_write -> SSEG_SEC_TENS:write_n
	wire  [31:0] mm_interconnect_0_sseg_sec_tens_s1_writedata;                 // mm_interconnect_0:SSEG_SEC_TENS_s1_writedata -> SSEG_SEC_TENS:writedata
	wire         mm_interconnect_0_sseg_hour_tens_s1_chipselect;               // mm_interconnect_0:SSEG_HOUR_TENS_s1_chipselect -> SSEG_HOUR_TENS:chipselect
	wire  [31:0] mm_interconnect_0_sseg_hour_tens_s1_readdata;                 // SSEG_HOUR_TENS:readdata -> mm_interconnect_0:SSEG_HOUR_TENS_s1_readdata
	wire   [1:0] mm_interconnect_0_sseg_hour_tens_s1_address;                  // mm_interconnect_0:SSEG_HOUR_TENS_s1_address -> SSEG_HOUR_TENS:address
	wire         mm_interconnect_0_sseg_hour_tens_s1_write;                    // mm_interconnect_0:SSEG_HOUR_TENS_s1_write -> SSEG_HOUR_TENS:write_n
	wire  [31:0] mm_interconnect_0_sseg_hour_tens_s1_writedata;                // mm_interconnect_0:SSEG_HOUR_TENS_s1_writedata -> SSEG_HOUR_TENS:writedata
	wire  [31:0] mm_interconnect_0_switch_s1_readdata;                         // SWITCH:readdata -> mm_interconnect_0:SWITCH_s1_readdata
	wire   [1:0] mm_interconnect_0_switch_s1_address;                          // mm_interconnect_0:SWITCH_s1_address -> SWITCH:address
	wire         mm_interconnect_0_buzzer_s1_chipselect;                       // mm_interconnect_0:BUZZER_s1_chipselect -> BUZZER:chipselect
	wire  [31:0] mm_interconnect_0_buzzer_s1_readdata;                         // BUZZER:readdata -> mm_interconnect_0:BUZZER_s1_readdata
	wire   [1:0] mm_interconnect_0_buzzer_s1_address;                          // mm_interconnect_0:BUZZER_s1_address -> BUZZER:address
	wire         mm_interconnect_0_buzzer_s1_write;                            // mm_interconnect_0:BUZZER_s1_write -> BUZZER:write_n
	wire  [31:0] mm_interconnect_0_buzzer_s1_writedata;                        // mm_interconnect_0:BUZZER_s1_writedata -> BUZZER:writedata
	wire         irq_mapper_receiver0_irq;                                     // DEBUG:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] timerwithclock_irq_irq;                                       // irq_mapper:sender_irq -> TimerWithClock:irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [BUTTONS:reset_n, BUZZER:reset_n, DEBUG:rst_n, LEDS:reset_n, SSEG_HOUR_TENS:reset_n, SSEG_HOUR_UNITS:reset_n, SSEG_MINS_TENS:reset_n, SSEG_MIN_UNITS:reset_n, SSEG_SEC_TENS:reset_n, SSEG_SEC_UNITS:reset_n, SWITCH:reset_n, TIMER:reset_n, TimerWithClock:reset_n, irq_mapper:reset, mm_interconnect_0:TimerWithClock_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [TimerWithClock:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                           // rst_controller_001:reset_out -> [SRAM:reset, mm_interconnect_0:SRAM_reset1_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                       // rst_controller_001:reset_req -> SRAM:reset_req

	TimerWithClock_BUTTONS buttons (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_buttons_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_buttons_s1_readdata), //                    .readdata
		.in_port  (buttons_export)                         // external_connection.export
	);

	TimerWithClock_BUZZER buzzer (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_buzzer_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_buzzer_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_buzzer_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_buzzer_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_buzzer_s1_readdata),   //                    .readdata
		.out_port   (buzzer_export)                           // external_connection.export
	);

	TimerWithClock_DEBUG debug (
		.clk            (clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_debug_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_debug_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_debug_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                               //               irq.irq
	);

	TimerWithClock_LEDS leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	TimerWithClock_SRAM sram (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_sram_s1_address),      //     s1.address
		.clken      (mm_interconnect_0_sram_s1_clken),        //       .clken
		.chipselect (mm_interconnect_0_sram_s1_chipselect),   //       .chipselect
		.write      (mm_interconnect_0_sram_s1_write),        //       .write
		.readdata   (mm_interconnect_0_sram_s1_readdata),     //       .readdata
		.writedata  (mm_interconnect_0_sram_s1_writedata),    //       .writedata
		.byteenable (mm_interconnect_0_sram_s1_byteenable),   //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	TimerWithClock_SSEG_HOUR_TENS sseg_hour_tens (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_sseg_hour_tens_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sseg_hour_tens_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sseg_hour_tens_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sseg_hour_tens_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sseg_hour_tens_s1_readdata),   //                    .readdata
		.out_port   (sseg_hour_tens_export)                           // external_connection.export
	);

	TimerWithClock_SSEG_HOUR_TENS sseg_hour_units (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_sseg_hour_units_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sseg_hour_units_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sseg_hour_units_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sseg_hour_units_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sseg_hour_units_s1_readdata),   //                    .readdata
		.out_port   (sseg_hour_units_export)                           // external_connection.export
	);

	TimerWithClock_SSEG_HOUR_TENS sseg_mins_tens (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_sseg_mins_tens_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sseg_mins_tens_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sseg_mins_tens_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sseg_mins_tens_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sseg_mins_tens_s1_readdata),   //                    .readdata
		.out_port   (sseg_mins_tens_export)                           // external_connection.export
	);

	TimerWithClock_SSEG_HOUR_TENS sseg_min_units (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_sseg_min_units_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sseg_min_units_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sseg_min_units_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sseg_min_units_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sseg_min_units_s1_readdata),   //                    .readdata
		.out_port   (sseg_min_units_export)                           // external_connection.export
	);

	TimerWithClock_SSEG_HOUR_TENS sseg_sec_tens (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_sseg_sec_tens_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sseg_sec_tens_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sseg_sec_tens_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sseg_sec_tens_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sseg_sec_tens_s1_readdata),   //                    .readdata
		.out_port   (sseg_sec_tens_export)                           // external_connection.export
	);

	TimerWithClock_SSEG_HOUR_TENS sseg_sec_units (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_sseg_sec_units_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sseg_sec_units_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sseg_sec_units_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sseg_sec_units_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sseg_sec_units_s1_readdata),   //                    .readdata
		.out_port   (sseg_sec_units_export)                           // external_connection.export
	);

	TimerWithClock_SWITCH switch (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_switch_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switch_s1_readdata), //                    .readdata
		.in_port  (switch_export)                         // external_connection.export
	);

	TimerWithClock_TIMER timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        ()                                       //   irq.irq
	);

	TimerWithClock_TimerWithClock timerwithclock (
		.clk                                 (clk_clk),                                                      //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                              //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                           (timerwithclock_data_master_address),                           //               data_master.address
		.d_byteenable                        (timerwithclock_data_master_byteenable),                        //                          .byteenable
		.d_read                              (timerwithclock_data_master_read),                              //                          .read
		.d_readdata                          (timerwithclock_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (timerwithclock_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (timerwithclock_data_master_write),                             //                          .write
		.d_writedata                         (timerwithclock_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (timerwithclock_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (timerwithclock_instruction_master_address),                    //        instruction_master.address
		.i_read                              (timerwithclock_instruction_master_read),                       //                          .read
		.i_readdata                          (timerwithclock_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (timerwithclock_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (timerwithclock_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (timerwithclock_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_timerwithclock_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_timerwithclock_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_timerwithclock_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_timerwithclock_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_timerwithclock_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_timerwithclock_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_timerwithclock_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_timerwithclock_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                              // custom_instruction_master.readra
	);

	TimerWithClock_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                      //                                  clk_0_clk.clk
		.SRAM_reset1_reset_bridge_in_reset_reset          (rst_controller_001_reset_out_reset),                           //          SRAM_reset1_reset_bridge_in_reset.reset
		.TimerWithClock_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // TimerWithClock_reset_reset_bridge_in_reset.reset
		.TimerWithClock_data_master_address               (timerwithclock_data_master_address),                           //                 TimerWithClock_data_master.address
		.TimerWithClock_data_master_waitrequest           (timerwithclock_data_master_waitrequest),                       //                                           .waitrequest
		.TimerWithClock_data_master_byteenable            (timerwithclock_data_master_byteenable),                        //                                           .byteenable
		.TimerWithClock_data_master_read                  (timerwithclock_data_master_read),                              //                                           .read
		.TimerWithClock_data_master_readdata              (timerwithclock_data_master_readdata),                          //                                           .readdata
		.TimerWithClock_data_master_write                 (timerwithclock_data_master_write),                             //                                           .write
		.TimerWithClock_data_master_writedata             (timerwithclock_data_master_writedata),                         //                                           .writedata
		.TimerWithClock_data_master_debugaccess           (timerwithclock_data_master_debugaccess),                       //                                           .debugaccess
		.TimerWithClock_instruction_master_address        (timerwithclock_instruction_master_address),                    //          TimerWithClock_instruction_master.address
		.TimerWithClock_instruction_master_waitrequest    (timerwithclock_instruction_master_waitrequest),                //                                           .waitrequest
		.TimerWithClock_instruction_master_read           (timerwithclock_instruction_master_read),                       //                                           .read
		.TimerWithClock_instruction_master_readdata       (timerwithclock_instruction_master_readdata),                   //                                           .readdata
		.BUTTONS_s1_address                               (mm_interconnect_0_buttons_s1_address),                         //                                 BUTTONS_s1.address
		.BUTTONS_s1_readdata                              (mm_interconnect_0_buttons_s1_readdata),                        //                                           .readdata
		.BUZZER_s1_address                                (mm_interconnect_0_buzzer_s1_address),                          //                                  BUZZER_s1.address
		.BUZZER_s1_write                                  (mm_interconnect_0_buzzer_s1_write),                            //                                           .write
		.BUZZER_s1_readdata                               (mm_interconnect_0_buzzer_s1_readdata),                         //                                           .readdata
		.BUZZER_s1_writedata                              (mm_interconnect_0_buzzer_s1_writedata),                        //                                           .writedata
		.BUZZER_s1_chipselect                             (mm_interconnect_0_buzzer_s1_chipselect),                       //                                           .chipselect
		.DEBUG_avalon_jtag_slave_address                  (mm_interconnect_0_debug_avalon_jtag_slave_address),            //                    DEBUG_avalon_jtag_slave.address
		.DEBUG_avalon_jtag_slave_write                    (mm_interconnect_0_debug_avalon_jtag_slave_write),              //                                           .write
		.DEBUG_avalon_jtag_slave_read                     (mm_interconnect_0_debug_avalon_jtag_slave_read),               //                                           .read
		.DEBUG_avalon_jtag_slave_readdata                 (mm_interconnect_0_debug_avalon_jtag_slave_readdata),           //                                           .readdata
		.DEBUG_avalon_jtag_slave_writedata                (mm_interconnect_0_debug_avalon_jtag_slave_writedata),          //                                           .writedata
		.DEBUG_avalon_jtag_slave_waitrequest              (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest),        //                                           .waitrequest
		.DEBUG_avalon_jtag_slave_chipselect               (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),         //                                           .chipselect
		.LEDS_s1_address                                  (mm_interconnect_0_leds_s1_address),                            //                                    LEDS_s1.address
		.LEDS_s1_write                                    (mm_interconnect_0_leds_s1_write),                              //                                           .write
		.LEDS_s1_readdata                                 (mm_interconnect_0_leds_s1_readdata),                           //                                           .readdata
		.LEDS_s1_writedata                                (mm_interconnect_0_leds_s1_writedata),                          //                                           .writedata
		.LEDS_s1_chipselect                               (mm_interconnect_0_leds_s1_chipselect),                         //                                           .chipselect
		.SRAM_s1_address                                  (mm_interconnect_0_sram_s1_address),                            //                                    SRAM_s1.address
		.SRAM_s1_write                                    (mm_interconnect_0_sram_s1_write),                              //                                           .write
		.SRAM_s1_readdata                                 (mm_interconnect_0_sram_s1_readdata),                           //                                           .readdata
		.SRAM_s1_writedata                                (mm_interconnect_0_sram_s1_writedata),                          //                                           .writedata
		.SRAM_s1_byteenable                               (mm_interconnect_0_sram_s1_byteenable),                         //                                           .byteenable
		.SRAM_s1_chipselect                               (mm_interconnect_0_sram_s1_chipselect),                         //                                           .chipselect
		.SRAM_s1_clken                                    (mm_interconnect_0_sram_s1_clken),                              //                                           .clken
		.SSEG_HOUR_TENS_s1_address                        (mm_interconnect_0_sseg_hour_tens_s1_address),                  //                          SSEG_HOUR_TENS_s1.address
		.SSEG_HOUR_TENS_s1_write                          (mm_interconnect_0_sseg_hour_tens_s1_write),                    //                                           .write
		.SSEG_HOUR_TENS_s1_readdata                       (mm_interconnect_0_sseg_hour_tens_s1_readdata),                 //                                           .readdata
		.SSEG_HOUR_TENS_s1_writedata                      (mm_interconnect_0_sseg_hour_tens_s1_writedata),                //                                           .writedata
		.SSEG_HOUR_TENS_s1_chipselect                     (mm_interconnect_0_sseg_hour_tens_s1_chipselect),               //                                           .chipselect
		.SSEG_HOUR_UNITS_s1_address                       (mm_interconnect_0_sseg_hour_units_s1_address),                 //                         SSEG_HOUR_UNITS_s1.address
		.SSEG_HOUR_UNITS_s1_write                         (mm_interconnect_0_sseg_hour_units_s1_write),                   //                                           .write
		.SSEG_HOUR_UNITS_s1_readdata                      (mm_interconnect_0_sseg_hour_units_s1_readdata),                //                                           .readdata
		.SSEG_HOUR_UNITS_s1_writedata                     (mm_interconnect_0_sseg_hour_units_s1_writedata),               //                                           .writedata
		.SSEG_HOUR_UNITS_s1_chipselect                    (mm_interconnect_0_sseg_hour_units_s1_chipselect),              //                                           .chipselect
		.SSEG_MIN_UNITS_s1_address                        (mm_interconnect_0_sseg_min_units_s1_address),                  //                          SSEG_MIN_UNITS_s1.address
		.SSEG_MIN_UNITS_s1_write                          (mm_interconnect_0_sseg_min_units_s1_write),                    //                                           .write
		.SSEG_MIN_UNITS_s1_readdata                       (mm_interconnect_0_sseg_min_units_s1_readdata),                 //                                           .readdata
		.SSEG_MIN_UNITS_s1_writedata                      (mm_interconnect_0_sseg_min_units_s1_writedata),                //                                           .writedata
		.SSEG_MIN_UNITS_s1_chipselect                     (mm_interconnect_0_sseg_min_units_s1_chipselect),               //                                           .chipselect
		.SSEG_MINS_TENS_s1_address                        (mm_interconnect_0_sseg_mins_tens_s1_address),                  //                          SSEG_MINS_TENS_s1.address
		.SSEG_MINS_TENS_s1_write                          (mm_interconnect_0_sseg_mins_tens_s1_write),                    //                                           .write
		.SSEG_MINS_TENS_s1_readdata                       (mm_interconnect_0_sseg_mins_tens_s1_readdata),                 //                                           .readdata
		.SSEG_MINS_TENS_s1_writedata                      (mm_interconnect_0_sseg_mins_tens_s1_writedata),                //                                           .writedata
		.SSEG_MINS_TENS_s1_chipselect                     (mm_interconnect_0_sseg_mins_tens_s1_chipselect),               //                                           .chipselect
		.SSEG_SEC_TENS_s1_address                         (mm_interconnect_0_sseg_sec_tens_s1_address),                   //                           SSEG_SEC_TENS_s1.address
		.SSEG_SEC_TENS_s1_write                           (mm_interconnect_0_sseg_sec_tens_s1_write),                     //                                           .write
		.SSEG_SEC_TENS_s1_readdata                        (mm_interconnect_0_sseg_sec_tens_s1_readdata),                  //                                           .readdata
		.SSEG_SEC_TENS_s1_writedata                       (mm_interconnect_0_sseg_sec_tens_s1_writedata),                 //                                           .writedata
		.SSEG_SEC_TENS_s1_chipselect                      (mm_interconnect_0_sseg_sec_tens_s1_chipselect),                //                                           .chipselect
		.SSEG_SEC_UNITS_s1_address                        (mm_interconnect_0_sseg_sec_units_s1_address),                  //                          SSEG_SEC_UNITS_s1.address
		.SSEG_SEC_UNITS_s1_write                          (mm_interconnect_0_sseg_sec_units_s1_write),                    //                                           .write
		.SSEG_SEC_UNITS_s1_readdata                       (mm_interconnect_0_sseg_sec_units_s1_readdata),                 //                                           .readdata
		.SSEG_SEC_UNITS_s1_writedata                      (mm_interconnect_0_sseg_sec_units_s1_writedata),                //                                           .writedata
		.SSEG_SEC_UNITS_s1_chipselect                     (mm_interconnect_0_sseg_sec_units_s1_chipselect),               //                                           .chipselect
		.SWITCH_s1_address                                (mm_interconnect_0_switch_s1_address),                          //                                  SWITCH_s1.address
		.SWITCH_s1_readdata                               (mm_interconnect_0_switch_s1_readdata),                         //                                           .readdata
		.TIMER_s1_address                                 (mm_interconnect_0_timer_s1_address),                           //                                   TIMER_s1.address
		.TIMER_s1_write                                   (mm_interconnect_0_timer_s1_write),                             //                                           .write
		.TIMER_s1_readdata                                (mm_interconnect_0_timer_s1_readdata),                          //                                           .readdata
		.TIMER_s1_writedata                               (mm_interconnect_0_timer_s1_writedata),                         //                                           .writedata
		.TIMER_s1_chipselect                              (mm_interconnect_0_timer_s1_chipselect),                        //                                           .chipselect
		.TimerWithClock_debug_mem_slave_address           (mm_interconnect_0_timerwithclock_debug_mem_slave_address),     //             TimerWithClock_debug_mem_slave.address
		.TimerWithClock_debug_mem_slave_write             (mm_interconnect_0_timerwithclock_debug_mem_slave_write),       //                                           .write
		.TimerWithClock_debug_mem_slave_read              (mm_interconnect_0_timerwithclock_debug_mem_slave_read),        //                                           .read
		.TimerWithClock_debug_mem_slave_readdata          (mm_interconnect_0_timerwithclock_debug_mem_slave_readdata),    //                                           .readdata
		.TimerWithClock_debug_mem_slave_writedata         (mm_interconnect_0_timerwithclock_debug_mem_slave_writedata),   //                                           .writedata
		.TimerWithClock_debug_mem_slave_byteenable        (mm_interconnect_0_timerwithclock_debug_mem_slave_byteenable),  //                                           .byteenable
		.TimerWithClock_debug_mem_slave_waitrequest       (mm_interconnect_0_timerwithclock_debug_mem_slave_waitrequest), //                                           .waitrequest
		.TimerWithClock_debug_mem_slave_debugaccess       (mm_interconnect_0_timerwithclock_debug_mem_slave_debugaccess)  //                                           .debugaccess
	);

	TimerWithClock_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (timerwithclock_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (timerwithclock_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),           // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),       //          .reset_req
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_in1      (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_in2      (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (timerwithclock_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                                  //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),       // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req),   //          .reset_req
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_in1      (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_in2      (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

endmodule
